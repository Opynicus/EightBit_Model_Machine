LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_ARITH.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY PC IS --程序计数器
PORT( 
 IPC,CLK,CLR:IN STD_LOGIC; 
 PC_out:OUT STD_LOGIC_VECTOR(3 DOWNTO 0) 
 ); 
END PC; 
ARCHITECTURE PC_arch OF PC IS 
SIGNAL tmp_out: STD_LOGIC_VECTOR(3 DOWNTO 0); 
BEGIN 
 PROCESS(CLK,CLR,IPC) 
 BEGIN 
 IF (CLR='0') THEN 
	tmp_out<= "0000"; 
 ELSIF (CLK'EVENT AND CLK='1') THEN 
	IF (IPC='1') THEN 
		tmp_out<= tmp_out+1; --PC+1 
	END IF; 
 END IF; 
 END PROCESS; 
 PC_out<= tmp_out; 
END PC_arch;