LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_ARITH.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 

ENTITY RAM IS 
 PORT( 
	DIN:IN STD_LOGIC_VECTOR(7 DOWNTO 0); --输入的内存内容
	DOUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0); --输出的是选中地址中相应的内容
	ADDR:IN STD_LOGIC_VECTOR(3 DOWNTO 0) ); --输入信号为地址信息
END RAM; 

ARCHITECTURE A OF RAM IS 
TYPE MEMORY IS ARRAY(0 TO 9) OF STD_LOGIC_VECTOR(7 DOWNTO 0); 
BEGIN 
	PROCESS(ADDR) 
	VARIABLE MEM: MEMORY; 
	BEGIN 
	MEM(0):="11000001";	--LD A,2H;
	MEM(1):="00000010";
	MEM(2):="11000010";	--ADD A,DH		
	MEM(3):="00001101";	
	MEM(4):="11000011";	--SUB A,4H;
	MEM(5):="00000101";
	MEM(6):="11000100";	--AND A,4H;
	MEM(7):="00000101";
	MEM(8):="11000101";	--SHL A,1;
	MEM(9):="11000000"; --停机
	DOUT <= MEM(CONV_INTEGER(ADDR(3 DOWNTO 0))); 
	END PROCESS; 
END A;