LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_ARITH.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 

ENTITY RAM IS 
 PORT( 
	WR,CS:IN STD_LOGIC; --WR片选信号, CS读写控制端
	DATA_IN:IN STD_LOGIC_VECTOR(7 DOWNTO 0); --输入的内存内容
	DATA_OUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0); --输出的是选中地址中相应的内容
	Address:IN STD_LOGIC_VECTOR(5 DOWNTO 0) ); --输入信号为地址信息
END RAM; 

ARCHITECTURE RAM_arch OF RAM IS 
TYPE MEMORY IS ARRAY(0 TO 34) OF STD_LOGIC_VECTOR(7 DOWNTO 0); 
BEGIN 
	PROCESS(CS,WR,Address) 
	VARIABLE MEM: MEMORY; 
	BEGIN 
	MEM(0):="00111110";	--LD A,6;
	MEM(1):="00000110";
	MEM(2):="11000110";	--ADD A,7		
	MEM(3):="00000111";	
	MEM(4):="00111110";	--LD A,7;
	MEM(5):="00000111";
	MEM(6):="00110011";	--SUB A,6
	MEM(7):="00000110";
	MEM(8):="00111110";	--LD A,6;
	MEM(9):="00000110";
	MEM(10):="01110001"; --AND A,7
	MEM(11):="00000111";
	MEM(12):="10110110"; --OR A,7
	MEM(13):="00000111";
	MEM(14):="00111110";	--LD A,7;
	MEM(15):="00000111";
	MEM(16):="10110110"; --OR A,8
	MEM(17):="00001000";
	MEM(18):="00111110";--LD A,8;
	MEM(19):="00001000";
	MEM(20):="01110110"; --XOR A,1
	MEM(21):="00000001";
	MEM(22):="00111110";--LD A,4;
	MEM(23):="00000100";
	MEM(24):="11000001";--NOT A
	MEM(25):="00111110";--LD A,4;
	MEM(26):="00000100";
	MEM(27):="11000010"; --NEG A
	MEM(28):="00111110";	--LD A,3;
	MEM(29):="00000011";
	MEM(30):="11000011"; --SHL
	MEM(31):="00111110";	--LD A,3;
	MEM(32):="00000011";
	MEM(33):="11000100"; --SHR
	MEM(34):="11000101"; --停机
	IF (CS='0') THEN 
		IF (WR='0') THEN 
			MEM(CONV_INTEGER(Address(5 DOWNTO 0))):=DATA_IN; 
		ELSIF(WR='1') THEN 
			DATA_OUT <= MEM(CONV_INTEGER(Address(5 DOWNTO 0))); 
		END IF; 
	END IF; 
	END PROCESS; 
END RAM_arch;