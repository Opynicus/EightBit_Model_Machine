LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 

ENTITY ACC IS --累加器模块
PORT( 
	DATA_IN:IN STD_LOGIC_VECTOR(7 DOWNTO 0); --输入
	IA:IN STD_LOGIC; --输入控制信号
	EA:IN STD_LOGIC; --输出控制信号
	CLK:IN STD_LOGIC; 
	DATA_OUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0) ); --输出
END ACC; 

ARCHITECTURE ACC_arch OF ACC IS 
SIGNAL REGQ : STD_LOGIC_VECTOR(7 DOWNTO 0); --中间信号
BEGIN 
	PROCESS(CLK,IA,EA,DATA_IN) 
	BEGIN 
	IF(CLK'EVENT AND CLK='1') THEN 
		IF(IA='0') THEN 
			REGQ<=DATA_IN; 
		END IF; 
	END IF; 
	END PROCESS; 
	DATA_OUT<=REGQ WHEN EA='0' ELSE "ZZZZZZZZ"; 
END ACC_arch;